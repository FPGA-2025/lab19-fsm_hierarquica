module sistema(
    input clk,
    input reset,
    input vai_manual,
    input vai_auto,
    input ligar_caldeira,
    output caldeira
);

// Insira seu código aqui

endmodule